
//Verilog file of module addSub


`timescale 1 ns / 1ns

module addSub_net(A,
B,
sel,
Result);
	input sel;
input [0:7]A;
input [0:7]B;
output [0:8]Result;
wire
addSub_wire_1,
addSub_wire_2,
addSub_wire_3,
addSub_wire_4,
addSub_wire_5,
addSub_wire_6,
addSub_wire_7,
addSub_wire_8,
addSub_wire_9,
addSub_wire_10,
addSub_wire_11,
addSub_wire_12,
addSub_wire_13,
addSub_wire_14,
addSub_wire_15,
addSub_wire_16,
addSub_wire_17,
addSub_wire_18,
addSub_wire_19,
addSub_wire_20,
addSub_wire_21,
addSub_wire_22,
addSub_wire_23,
addSub_wire_24,
addSub_wire_25,
addSub_wire_26,
addSub_wire_27,
addSub_wire_28,
addSub_wire_29,
addSub_wire_30,
addSub_wire_31,
addSub_wire_32,
addSub_wire_33,
addSub_wire_34,
addSub_wire_35,
addSub_wire_36,
addSub_wire_37,
addSub_wire_38,
addSub_wire_39,
addSub_wire_40,
addSub_wire_41,
addSub_wire_42,
addSub_wire_43,
addSub_wire_44,
addSub_wire_45,
addSub_wire_46,
addSub_wire_47,
addSub_wire_48,
addSub_wire_49,
addSub_wire_50,
addSub_wire_51,
addSub_wire_52,
addSub_wire_53,
addSub_wire_54,
addSub_wire_55,
addSub_wire_56,
addSub_wire_57,
addSub_wire_58,
addSub_wire_59,
addSub_wire_60,
addSub_wire_61,
addSub_wire_62,
addSub_wire_63,
addSub_wire_64,
addSub_wire_65,
addSub_wire_66,
addSub_wire_67,
addSub_wire_68,
addSub_wire_69,
addSub_wire_70,
addSub_wire_71,
addSub_wire_72,
addSub_wire_73,
addSub_wire_74,
addSub_wire_75,
addSub_wire_76,
addSub_wire_77,
addSub_wire_78,
addSub_wire_79,
addSub_wire_80,
addSub_wire_81,
addSub_wire_82,
addSub_wire_83,
addSub_wire_84,
addSub_wire_85,
addSub_wire_86,
addSub_wire_87,
addSub_wire_88,
addSub_wire_89,
addSub_wire_90,
addSub_wire_91,
addSub_wire_92,
addSub_wire_93,
addSub_wire_94,
addSub_wire_95,
addSub_wire_96,
addSub_wire_97,
addSub_wire_98,
addSub_wire_99,
addSub_wire_100,
addSub_wire_101,
addSub_wire_102,
addSub_wire_103,
addSub_wire_104,
addSub_wire_105,
addSub_wire_106,
addSub_wire_107,
addSub_wire_108,
addSub_wire_109,
addSub_wire_110,
addSub_wire_111,
addSub_wire_112,
addSub_wire_113,
addSub_wire_114,
addSub_wire_115,
addSub_wire_116,
addSub_wire_117,
addSub_wire_118,
addSub_wire_119,
addSub_wire_120,
addSub_wire_121,
addSub_wire_122,
addSub_wire_123,
addSub_wire_124,
addSub_wire_125,
addSub_wire_126,
addSub_wire_127,
addSub_wire_128,
addSub_wire_129,
addSub_wire_130,
addSub_wire_131,
addSub_wire_132,
addSub_wire_133,
addSub_wire_134,
addSub_wire_135,
addSub_wire_136,
addSub_wire_137,
addSub_wire_138,
addSub_wire_139,
addSub_wire_140,
addSub_wire_141,
addSub_wire_142,
addSub_wire_143,
addSub_wire_144,
addSub_wire_145,
addSub_wire_146,
addSub_wire_147,
addSub_wire_148,
addSub_wire_149,
addSub_wire_150,
addSub_wire_151,
addSub_wire_152,
addSub_wire_153,
addSub_wire_154,
addSub_wire_3_0,
addSub_wire_3_1,
addSub_wire_3_2,
addSub_wire_3_3,
addSub_wire_37_0,
addSub_wire_37_1,
addSub_wire_37_2,
addSub_wire_37_3,
addSub_wire_32_0,
addSub_wire_32_1,
addSub_wire_32_2,
addSub_wire_32_3,
addSub_wire_27_0,
addSub_wire_27_1,
addSub_wire_27_2,
addSub_wire_27_3,
addSub_wire_22_0,
addSub_wire_22_1,
addSub_wire_22_2,
addSub_wire_22_3,
addSub_wire_17_0,
addSub_wire_17_1,
addSub_wire_17_2,
addSub_wire_17_3,
addSub_wire_12_0,
addSub_wire_12_1,
addSub_wire_12_2,
addSub_wire_12_3,
addSub_wire_7_0,
addSub_wire_7_1,
addSub_wire_7_2,
addSub_wire_7_3,
addSub_wire_60_0,
addSub_wire_60_1,
addSub_wire_60_2,
addSub_wire_36_0,
addSub_wire_36_1,
addSub_wire_36_2,
addSub_wire_2_0,
addSub_wire_2_1,
addSub_wire_2_2,
addSub_wire_2_3,
addSub_wire_38_0,
addSub_wire_38_1,
addSub_wire_38_2,
addSub_wire_38_3,
addSub_wire_38_4,
addSub_wire_38_5,
addSub_wire_33_0,
addSub_wire_33_1,
addSub_wire_33_2,
addSub_wire_33_3,
addSub_wire_33_4,
addSub_wire_33_5,
addSub_wire_28_0,
addSub_wire_28_1,
addSub_wire_28_2,
addSub_wire_28_3,
addSub_wire_28_4,
addSub_wire_28_5,
addSub_wire_23_0,
addSub_wire_23_1,
addSub_wire_23_2,
addSub_wire_23_3,
addSub_wire_23_4,
addSub_wire_23_5,
addSub_wire_18_0,
addSub_wire_18_1,
addSub_wire_18_2,
addSub_wire_18_3,
addSub_wire_18_4,
addSub_wire_18_5,
addSub_wire_13_0,
addSub_wire_13_1,
addSub_wire_13_2,
addSub_wire_13_3,
addSub_wire_13_4,
addSub_wire_13_5,
addSub_wire_8_0,
addSub_wire_8_1,
addSub_wire_8_2,
addSub_wire_8_3,
addSub_wire_8_4,
addSub_wire_8_5,
addSub_wire_31_0,
addSub_wire_31_1,
addSub_wire_31_2,
addSub_wire_26_0,
addSub_wire_26_1,
addSub_wire_26_2,
addSub_wire_21_0,
addSub_wire_21_1,
addSub_wire_21_2,
addSub_wire_16_0,
addSub_wire_16_1,
addSub_wire_16_2,
addSub_wire_11_0,
addSub_wire_11_1,
addSub_wire_11_2,
addSub_wire_6_0,
addSub_wire_6_1,
addSub_wire_6_2,
addSub_wire_57_0,
addSub_wire_57_1,
addSub_wire_57_2,
addSub_wire_54_0,
addSub_wire_54_1,
addSub_wire_54_2,
addSub_wire_51_0,
addSub_wire_51_1,
addSub_wire_51_2,
addSub_wire_48_0,
addSub_wire_48_1,
addSub_wire_48_2,
addSub_wire_45_0,
addSub_wire_45_1,
addSub_wire_45_2,
addSub_wire_42_0,
addSub_wire_42_1,
addSub_wire_42_2,
addSub_wire_121_0,
addSub_wire_121_1,
addSub_wire_121_2,
addSub_wire_121_3,
addSub_wire_121_4,
addSub_wire_121_5,
addSub_wire_121_6,
addSub_wire_121_7,
addSub_wire_121_8,
addSub_wire_121_9,
addSub_wire_121_10,
addSub_wire_121_11,
addSub_wire_121_12,
addSub_wire_121_13,
addSub_wire_121_14,
addSub_wire_121_15,
addSub_wire_121_16,
addSub_wire_121_17,
sel_net_0;

pin #(17) pin_0 ({sel, A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], B[0], B[1], B[2], B[3], B[4], B[5], B[6], B[7]}, {sel_net_0, A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, B_0, B_1, B_2, B_3, B_4, B_5, B_6, B_7});

pout #(9) pout_0 ({Result_0, Result_1, Result_2, Result_3, Result_4, Result_5, Result_6, Result_7, Result_8}, {Result[0], Result[1], Result[2], Result[3], Result[4], Result[5], Result[6], Result[7], Result[8]});

fanout_n #(4, 0, 0) FANOUT_1 (addSub_wire_3, {addSub_wire_3_0, addSub_wire_3_1, addSub_wire_3_2, addSub_wire_3_3});
fanout_n #(4, 0, 0) FANOUT_2 (addSub_wire_37, {addSub_wire_37_0, addSub_wire_37_1, addSub_wire_37_2, addSub_wire_37_3});
fanout_n #(4, 0, 0) FANOUT_3 (addSub_wire_32, {addSub_wire_32_0, addSub_wire_32_1, addSub_wire_32_2, addSub_wire_32_3});
fanout_n #(4, 0, 0) FANOUT_4 (addSub_wire_27, {addSub_wire_27_0, addSub_wire_27_1, addSub_wire_27_2, addSub_wire_27_3});
fanout_n #(4, 0, 0) FANOUT_5 (addSub_wire_22, {addSub_wire_22_0, addSub_wire_22_1, addSub_wire_22_2, addSub_wire_22_3});
fanout_n #(4, 0, 0) FANOUT_6 (addSub_wire_17, {addSub_wire_17_0, addSub_wire_17_1, addSub_wire_17_2, addSub_wire_17_3});
fanout_n #(4, 0, 0) FANOUT_7 (addSub_wire_12, {addSub_wire_12_0, addSub_wire_12_1, addSub_wire_12_2, addSub_wire_12_3});
fanout_n #(4, 0, 0) FANOUT_8 (addSub_wire_7, {addSub_wire_7_0, addSub_wire_7_1, addSub_wire_7_2, addSub_wire_7_3});
fanout_n #(3, 0, 0) FANOUT_9 (addSub_wire_60, {addSub_wire_60_0, addSub_wire_60_1, addSub_wire_60_2});
fanout_n #(3, 0, 0) FANOUT_10 (addSub_wire_36, {addSub_wire_36_0, addSub_wire_36_1, addSub_wire_36_2});
fanout_n #(4, 0, 0) FANOUT_11 (addSub_wire_2, {addSub_wire_2_0, addSub_wire_2_1, addSub_wire_2_2, addSub_wire_2_3});
fanout_n #(6, 0, 0) FANOUT_12 (addSub_wire_38, {addSub_wire_38_0, addSub_wire_38_1, addSub_wire_38_2, addSub_wire_38_3, addSub_wire_38_4, addSub_wire_38_5});
fanout_n #(6, 0, 0) FANOUT_13 (addSub_wire_33, {addSub_wire_33_0, addSub_wire_33_1, addSub_wire_33_2, addSub_wire_33_3, addSub_wire_33_4, addSub_wire_33_5});
fanout_n #(6, 0, 0) FANOUT_14 (addSub_wire_28, {addSub_wire_28_0, addSub_wire_28_1, addSub_wire_28_2, addSub_wire_28_3, addSub_wire_28_4, addSub_wire_28_5});
fanout_n #(6, 0, 0) FANOUT_15 (addSub_wire_23, {addSub_wire_23_0, addSub_wire_23_1, addSub_wire_23_2, addSub_wire_23_3, addSub_wire_23_4, addSub_wire_23_5});
fanout_n #(6, 0, 0) FANOUT_16 (addSub_wire_18, {addSub_wire_18_0, addSub_wire_18_1, addSub_wire_18_2, addSub_wire_18_3, addSub_wire_18_4, addSub_wire_18_5});
fanout_n #(6, 0, 0) FANOUT_17 (addSub_wire_13, {addSub_wire_13_0, addSub_wire_13_1, addSub_wire_13_2, addSub_wire_13_3, addSub_wire_13_4, addSub_wire_13_5});
fanout_n #(6, 0, 0) FANOUT_18 (addSub_wire_8, {addSub_wire_8_0, addSub_wire_8_1, addSub_wire_8_2, addSub_wire_8_3, addSub_wire_8_4, addSub_wire_8_5});
fanout_n #(3, 0, 0) FANOUT_19 (addSub_wire_31, {addSub_wire_31_0, addSub_wire_31_1, addSub_wire_31_2});
fanout_n #(3, 0, 0) FANOUT_20 (addSub_wire_26, {addSub_wire_26_0, addSub_wire_26_1, addSub_wire_26_2});
fanout_n #(3, 0, 0) FANOUT_21 (addSub_wire_21, {addSub_wire_21_0, addSub_wire_21_1, addSub_wire_21_2});
fanout_n #(3, 0, 0) FANOUT_22 (addSub_wire_16, {addSub_wire_16_0, addSub_wire_16_1, addSub_wire_16_2});
fanout_n #(3, 0, 0) FANOUT_23 (addSub_wire_11, {addSub_wire_11_0, addSub_wire_11_1, addSub_wire_11_2});
fanout_n #(3, 0, 0) FANOUT_24 (addSub_wire_6, {addSub_wire_6_0, addSub_wire_6_1, addSub_wire_6_2});
fanout_n #(3, 0, 0) FANOUT_25 (addSub_wire_57, {addSub_wire_57_0, addSub_wire_57_1, addSub_wire_57_2});
fanout_n #(3, 0, 0) FANOUT_26 (addSub_wire_54, {addSub_wire_54_0, addSub_wire_54_1, addSub_wire_54_2});
fanout_n #(3, 0, 0) FANOUT_27 (addSub_wire_51, {addSub_wire_51_0, addSub_wire_51_1, addSub_wire_51_2});
fanout_n #(3, 0, 0) FANOUT_28 (addSub_wire_48, {addSub_wire_48_0, addSub_wire_48_1, addSub_wire_48_2});
fanout_n #(3, 0, 0) FANOUT_29 (addSub_wire_45, {addSub_wire_45_0, addSub_wire_45_1, addSub_wire_45_2});
fanout_n #(3, 0, 0) FANOUT_30 (addSub_wire_42, {addSub_wire_42_0, addSub_wire_42_1, addSub_wire_42_2});
fanout_n #(18, 0, 0) FANOUT_31 (addSub_wire_121, {addSub_wire_121_0, addSub_wire_121_1, addSub_wire_121_2, addSub_wire_121_3, addSub_wire_121_4, addSub_wire_121_5, addSub_wire_121_6, addSub_wire_121_7, addSub_wire_121_8, addSub_wire_121_9, addSub_wire_121_10, addSub_wire_121_11, addSub_wire_121_12, addSub_wire_121_13, addSub_wire_121_14, addSub_wire_121_15, addSub_wire_121_16, addSub_wire_121_17});


xor_n #(2, 0, 0) XOR_1 (addSub_wire_1, {addSub_wire_2_0, addSub_wire_3_0});
xor_n #(2, 0, 0) XOR_2 (addSub_wire_4, {addSub_wire_5, addSub_wire_6_0});
xor_n #(2, 0, 0) XOR_3 (addSub_wire_5, {addSub_wire_7_0, addSub_wire_8_0});
xor_n #(2, 0, 0) XOR_4 (addSub_wire_9, {addSub_wire_10, addSub_wire_11_0});
xor_n #(2, 0, 0) XOR_5 (addSub_wire_10, {addSub_wire_12_0, addSub_wire_13_0});
xor_n #(2, 0, 0) XOR_6 (addSub_wire_14, {addSub_wire_15, addSub_wire_16_0});
xor_n #(2, 0, 0) XOR_7 (addSub_wire_15, {addSub_wire_17_0, addSub_wire_18_0});
xor_n #(2, 0, 0) XOR_8 (addSub_wire_19, {addSub_wire_20, addSub_wire_21_0});
xor_n #(2, 0, 0) XOR_9 (addSub_wire_20, {addSub_wire_22_0, addSub_wire_23_0});
xor_n #(2, 0, 0) XOR_10 (addSub_wire_24, {addSub_wire_25, addSub_wire_26_0});
xor_n #(2, 0, 0) XOR_11 (addSub_wire_25, {addSub_wire_27_0, addSub_wire_28_0});
xor_n #(2, 0, 0) XOR_12 (addSub_wire_29, {addSub_wire_30, addSub_wire_31_0});
xor_n #(2, 0, 0) XOR_13 (addSub_wire_30, {addSub_wire_32_0, addSub_wire_33_0});
xor_n #(2, 0, 0) XOR_14 (addSub_wire_34, {addSub_wire_35, addSub_wire_36_0});
xor_n #(2, 0, 0) XOR_15 (addSub_wire_35, {addSub_wire_37_0, addSub_wire_38_0});
xnor_n #(2, 0, 0) XNOR_1 (addSub_wire_39, {addSub_wire_2_1, addSub_wire_3_1});
xor_n #(2, 0, 0) XOR_16 (addSub_wire_40, {addSub_wire_41, addSub_wire_42_0});
xnor_n #(2, 0, 0) XNOR_2 (addSub_wire_41, {addSub_wire_7_1, addSub_wire_8_1});
xor_n #(2, 0, 0) XOR_17 (addSub_wire_43, {addSub_wire_44, addSub_wire_45_0});
xnor_n #(2, 0, 0) XNOR_3 (addSub_wire_44, {addSub_wire_12_1, addSub_wire_13_1});
xor_n #(2, 0, 0) XOR_18 (addSub_wire_46, {addSub_wire_47, addSub_wire_48_0});
xnor_n #(2, 0, 0) XNOR_4 (addSub_wire_47, {addSub_wire_17_1, addSub_wire_18_1});
xor_n #(2, 0, 0) XOR_19 (addSub_wire_49, {addSub_wire_50, addSub_wire_51_0});
xnor_n #(2, 0, 0) XNOR_5 (addSub_wire_50, {addSub_wire_22_1, addSub_wire_23_1});
xor_n #(2, 0, 0) XOR_20 (addSub_wire_52, {addSub_wire_53, addSub_wire_54_0});
xnor_n #(2, 0, 0) XNOR_6 (addSub_wire_53, {addSub_wire_27_1, addSub_wire_28_1});
xor_n #(2, 0, 0) XOR_21 (addSub_wire_55, {addSub_wire_56, addSub_wire_57_0});
xnor_n #(2, 0, 0) XNOR_7 (addSub_wire_56, {addSub_wire_32_1, addSub_wire_33_1});
xor_n #(2, 0, 0) XOR_22 (addSub_wire_58, {addSub_wire_59, addSub_wire_60_0});
xnor_n #(2, 0, 0) XNOR_8 (addSub_wire_59, {addSub_wire_37_1, addSub_wire_38_1});
bufg #(0, 0) BUF_1 (addSub_wire_3, A_7);
bufg #(0, 0) BUF_2 (addSub_wire_37, A_6);
bufg #(0, 0) BUF_3 (addSub_wire_32, A_5);
bufg #(0, 0) BUF_4 (addSub_wire_27, A_4);
bufg #(0, 0) BUF_5 (addSub_wire_22, A_3);
bufg #(0, 0) BUF_6 (addSub_wire_17, A_2);
bufg #(0, 0) BUF_7 (addSub_wire_12, A_1);
bufg #(0, 0) BUF_8 (addSub_wire_7, A_0);
or_n #(2, 0, 0) OR_1 (addSub_wire_60, {addSub_wire_3_2, addSub_wire_61});
and_n #(2, 0, 0) AND_1 (addSub_wire_36, {addSub_wire_3_3, addSub_wire_2_2});
and_n #(2, 0, 0) AND_2 (addSub_wire_62, {addSub_wire_37_2, addSub_wire_63});
and_n #(2, 0, 0) AND_3 (addSub_wire_64, {addSub_wire_37_3, addSub_wire_65});
and_n #(2, 0, 0) AND_4 (addSub_wire_66, {addSub_wire_32_2, addSub_wire_67});
and_n #(2, 0, 0) AND_5 (addSub_wire_68, {addSub_wire_32_3, addSub_wire_69});
and_n #(2, 0, 0) AND_6 (addSub_wire_70, {addSub_wire_27_2, addSub_wire_71});
and_n #(2, 0, 0) AND_7 (addSub_wire_72, {addSub_wire_27_3, addSub_wire_73});
and_n #(2, 0, 0) AND_8 (addSub_wire_74, {addSub_wire_22_2, addSub_wire_75});
and_n #(2, 0, 0) AND_9 (addSub_wire_76, {addSub_wire_22_3, addSub_wire_77});
and_n #(2, 0, 0) AND_10 (addSub_wire_78, {addSub_wire_17_2, addSub_wire_79});
and_n #(2, 0, 0) AND_11 (addSub_wire_80, {addSub_wire_17_3, addSub_wire_81});
and_n #(2, 0, 0) AND_12 (addSub_wire_82, {addSub_wire_12_2, addSub_wire_83});
and_n #(2, 0, 0) AND_13 (addSub_wire_84, {addSub_wire_12_3, addSub_wire_85});
and_n #(2, 0, 0) AND_14 (addSub_wire_86, {addSub_wire_7_2, addSub_wire_87});
and_n #(2, 0, 0) AND_15 (addSub_wire_88, {addSub_wire_7_3, addSub_wire_89});
bufg #(0, 0) BUF_9 (addSub_wire_2, B_7);
bufg #(0, 0) BUF_10 (addSub_wire_38, B_6);
bufg #(0, 0) BUF_11 (addSub_wire_33, B_5);
bufg #(0, 0) BUF_12 (addSub_wire_28, B_4);
bufg #(0, 0) BUF_13 (addSub_wire_23, B_3);
bufg #(0, 0) BUF_14 (addSub_wire_18, B_2);
bufg #(0, 0) BUF_15 (addSub_wire_13, B_1);
bufg #(0, 0) BUF_16 (addSub_wire_8, B_0);
notg #(0, 0) NOT_1 (addSub_wire_61, addSub_wire_2_3);
notg #(0, 0) NOT_2 (addSub_wire_90, addSub_wire_38_2);
notg #(0, 0) NOT_3 (addSub_wire_91, addSub_wire_38_3);
and_n #(2, 0, 0) AND_16 (addSub_wire_92, {addSub_wire_38_4, addSub_wire_36_1});
or_n #(2, 0, 0) OR_2 (addSub_wire_65, {addSub_wire_38_5, addSub_wire_36_2});
notg #(0, 0) NOT_4 (addSub_wire_93, addSub_wire_33_2);
notg #(0, 0) NOT_5 (addSub_wire_94, addSub_wire_33_3);
and_n #(2, 0, 0) AND_17 (addSub_wire_95, {addSub_wire_33_4, addSub_wire_31_1});
or_n #(2, 0, 0) OR_3 (addSub_wire_69, {addSub_wire_33_5, addSub_wire_31_2});
notg #(0, 0) NOT_6 (addSub_wire_96, addSub_wire_28_2);
notg #(0, 0) NOT_7 (addSub_wire_97, addSub_wire_28_3);
and_n #(2, 0, 0) AND_18 (addSub_wire_98, {addSub_wire_28_4, addSub_wire_26_1});
or_n #(2, 0, 0) OR_4 (addSub_wire_73, {addSub_wire_28_5, addSub_wire_26_2});
notg #(0, 0) NOT_8 (addSub_wire_99, addSub_wire_23_2);
notg #(0, 0) NOT_9 (addSub_wire_100, addSub_wire_23_3);
and_n #(2, 0, 0) AND_19 (addSub_wire_101, {addSub_wire_23_4, addSub_wire_21_1});
or_n #(2, 0, 0) OR_5 (addSub_wire_77, {addSub_wire_23_5, addSub_wire_21_2});
notg #(0, 0) NOT_10 (addSub_wire_102, addSub_wire_18_2);
notg #(0, 0) NOT_11 (addSub_wire_103, addSub_wire_18_3);
and_n #(2, 0, 0) AND_20 (addSub_wire_104, {addSub_wire_18_4, addSub_wire_16_1});
or_n #(2, 0, 0) OR_6 (addSub_wire_81, {addSub_wire_18_5, addSub_wire_16_2});
notg #(0, 0) NOT_12 (addSub_wire_105, addSub_wire_13_2);
notg #(0, 0) NOT_13 (addSub_wire_106, addSub_wire_13_3);
and_n #(2, 0, 0) AND_21 (addSub_wire_107, {addSub_wire_13_4, addSub_wire_11_1});
or_n #(2, 0, 0) OR_7 (addSub_wire_85, {addSub_wire_13_5, addSub_wire_11_2});
notg #(0, 0) NOT_14 (addSub_wire_108, addSub_wire_8_2);
notg #(0, 0) NOT_15 (addSub_wire_109, addSub_wire_8_3);
and_n #(2, 0, 0) AND_22 (addSub_wire_110, {addSub_wire_8_4, addSub_wire_6_1});
or_n #(2, 0, 0) OR_8 (addSub_wire_89, {addSub_wire_8_5, addSub_wire_6_2});
or_n #(2, 0, 0) OR_9 (addSub_wire_31, {addSub_wire_92, addSub_wire_64});
or_n #(2, 0, 0) OR_10 (addSub_wire_26, {addSub_wire_95, addSub_wire_68});
or_n #(2, 0, 0) OR_11 (addSub_wire_21, {addSub_wire_98, addSub_wire_72});
or_n #(2, 0, 0) OR_12 (addSub_wire_16, {addSub_wire_101, addSub_wire_76});
or_n #(2, 0, 0) OR_13 (addSub_wire_11, {addSub_wire_104, addSub_wire_80});
or_n #(2, 0, 0) OR_14 (addSub_wire_6, {addSub_wire_107, addSub_wire_84});
or_n #(2, 0, 0) OR_15 (addSub_wire_63, {addSub_wire_60_1, addSub_wire_90});
and_n #(2, 0, 0) AND_23 (addSub_wire_111, {addSub_wire_60_2, addSub_wire_91});
or_n #(2, 0, 0) OR_16 (addSub_wire_57, {addSub_wire_111, addSub_wire_62});
or_n #(2, 0, 0) OR_17 (addSub_wire_67, {addSub_wire_57_1, addSub_wire_93});
and_n #(2, 0, 0) AND_24 (addSub_wire_112, {addSub_wire_57_2, addSub_wire_94});
or_n #(2, 0, 0) OR_18 (addSub_wire_54, {addSub_wire_112, addSub_wire_66});
or_n #(2, 0, 0) OR_19 (addSub_wire_71, {addSub_wire_54_1, addSub_wire_96});
and_n #(2, 0, 0) AND_25 (addSub_wire_113, {addSub_wire_54_2, addSub_wire_97});
or_n #(2, 0, 0) OR_20 (addSub_wire_51, {addSub_wire_113, addSub_wire_70});
or_n #(2, 0, 0) OR_21 (addSub_wire_75, {addSub_wire_51_1, addSub_wire_99});
and_n #(2, 0, 0) AND_26 (addSub_wire_114, {addSub_wire_51_2, addSub_wire_100});
or_n #(2, 0, 0) OR_22 (addSub_wire_48, {addSub_wire_114, addSub_wire_74});
or_n #(2, 0, 0) OR_23 (addSub_wire_79, {addSub_wire_48_1, addSub_wire_102});
and_n #(2, 0, 0) AND_27 (addSub_wire_115, {addSub_wire_48_2, addSub_wire_103});
or_n #(2, 0, 0) OR_24 (addSub_wire_45, {addSub_wire_115, addSub_wire_78});
or_n #(2, 0, 0) OR_25 (addSub_wire_83, {addSub_wire_45_1, addSub_wire_105});
and_n #(2, 0, 0) AND_28 (addSub_wire_116, {addSub_wire_45_2, addSub_wire_106});
or_n #(2, 0, 0) OR_26 (addSub_wire_42, {addSub_wire_116, addSub_wire_82});
or_n #(2, 0, 0) OR_27 (addSub_wire_87, {addSub_wire_42_1, addSub_wire_108});
and_n #(2, 0, 0) AND_29 (addSub_wire_117, {addSub_wire_42_2, addSub_wire_109});
or_n #(2, 0, 0) OR_28 (addSub_wire_118, {addSub_wire_117, addSub_wire_86});
bufg #(0, 0) BUF_17 (Result_8, addSub_wire_119);
and_n #(2, 0, 0) AND_30 (addSub_wire_120, {addSub_wire_1, addSub_wire_121_0});
or_n #(2, 0, 0) OR_29 (addSub_wire_119, {addSub_wire_120, addSub_wire_122});
nor_n #(2, 0, 0) NOR_1 (addSub_wire_122, {addSub_wire_121_1, addSub_wire_39});
bufg #(0, 0) BUF_18 (Result_7, addSub_wire_123);
and_n #(2, 0, 0) AND_31 (addSub_wire_124, {addSub_wire_34, addSub_wire_121_2});
or_n #(2, 0, 0) OR_30 (addSub_wire_123, {addSub_wire_124, addSub_wire_125});
notg #(0, 0) NOT_16 (addSub_wire_126, addSub_wire_121_3);
and_n #(2, 0, 0) AND_32 (addSub_wire_125, {addSub_wire_126, addSub_wire_58});
bufg #(0, 0) BUF_19 (Result_6, addSub_wire_127);
and_n #(2, 0, 0) AND_33 (addSub_wire_128, {addSub_wire_29, addSub_wire_121_4});
or_n #(2, 0, 0) OR_31 (addSub_wire_127, {addSub_wire_128, addSub_wire_129});
notg #(0, 0) NOT_17 (addSub_wire_130, addSub_wire_121_5);
and_n #(2, 0, 0) AND_34 (addSub_wire_129, {addSub_wire_130, addSub_wire_55});
bufg #(0, 0) BUF_20 (Result_5, addSub_wire_131);
and_n #(2, 0, 0) AND_35 (addSub_wire_132, {addSub_wire_24, addSub_wire_121_6});
or_n #(2, 0, 0) OR_32 (addSub_wire_131, {addSub_wire_132, addSub_wire_133});
notg #(0, 0) NOT_18 (addSub_wire_134, addSub_wire_121_7);
and_n #(2, 0, 0) AND_36 (addSub_wire_133, {addSub_wire_134, addSub_wire_52});
bufg #(0, 0) BUF_21 (Result_4, addSub_wire_135);
and_n #(2, 0, 0) AND_37 (addSub_wire_136, {addSub_wire_19, addSub_wire_121_8});
or_n #(2, 0, 0) OR_33 (addSub_wire_135, {addSub_wire_136, addSub_wire_137});
notg #(0, 0) NOT_19 (addSub_wire_138, addSub_wire_121_9);
and_n #(2, 0, 0) AND_38 (addSub_wire_137, {addSub_wire_138, addSub_wire_49});
bufg #(0, 0) BUF_22 (Result_3, addSub_wire_139);
and_n #(2, 0, 0) AND_39 (addSub_wire_140, {addSub_wire_14, addSub_wire_121_10});
or_n #(2, 0, 0) OR_34 (addSub_wire_139, {addSub_wire_140, addSub_wire_141});
notg #(0, 0) NOT_20 (addSub_wire_142, addSub_wire_121_11);
and_n #(2, 0, 0) AND_40 (addSub_wire_141, {addSub_wire_142, addSub_wire_46});
bufg #(0, 0) BUF_23 (Result_2, addSub_wire_143);
and_n #(2, 0, 0) AND_41 (addSub_wire_144, {addSub_wire_9, addSub_wire_121_12});
or_n #(2, 0, 0) OR_35 (addSub_wire_143, {addSub_wire_144, addSub_wire_145});
notg #(0, 0) NOT_21 (addSub_wire_146, addSub_wire_121_13);
and_n #(2, 0, 0) AND_42 (addSub_wire_145, {addSub_wire_146, addSub_wire_43});
bufg #(0, 0) BUF_24 (Result_1, addSub_wire_147);
and_n #(2, 0, 0) AND_43 (addSub_wire_148, {addSub_wire_4, addSub_wire_121_14});
or_n #(2, 0, 0) OR_36 (addSub_wire_147, {addSub_wire_148, addSub_wire_149});
notg #(0, 0) NOT_22 (addSub_wire_150, addSub_wire_121_15);
and_n #(2, 0, 0) AND_44 (addSub_wire_149, {addSub_wire_150, addSub_wire_40});
bufg #(0, 0) BUF_25 (Result_0, addSub_wire_151);
or_n #(2, 0, 0) OR_37 (addSub_wire_152, {addSub_wire_110, addSub_wire_88});
nor_n #(2, 0, 0) NOR_2 (addSub_wire_153, {addSub_wire_121_16, addSub_wire_118});
or_n #(2, 0, 0) OR_38 (addSub_wire_151, {addSub_wire_153, addSub_wire_154});
and_n #(2, 0, 0) AND_45 (addSub_wire_154, {addSub_wire_152, addSub_wire_121_17});
bufg #(0, 0) BUF_26 (addSub_wire_121, sel_net_0);

endmodule
